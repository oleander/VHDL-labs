linus@dhcp-076097.eduroam.chalmers.se.25605