linus@banan.olf.sgsnet.se.97665