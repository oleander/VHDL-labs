linus@dhcp-079070.eduroam.chalmers.se.42077