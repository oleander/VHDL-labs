linus@linus-oleanders-macbook.local.60830