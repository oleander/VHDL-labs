linus@linus-oleanders-macbook.local.61810