linus@linus-oleanders-macbook.local.61683