library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity mealy is
  port (clk, reset : in  std_logic;
        x          : in  std_logic_vector(1 downto 0);
        u          : out std_logic;
        q, qp      : out std_logic_vector(1 downto 0)
        );
end mealy;

end entity;  -- mealy

architecture arch of mealy is

begin

end architecture;  -- arch
