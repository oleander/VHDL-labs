linus@linus-oleanders-macbook.local.71406