linus@dhcp-075015.eduroam.chalmers.se.24144