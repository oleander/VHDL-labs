linus@linus-oleanders-macbook.local.15000