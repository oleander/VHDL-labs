linus@dhcp-078062.eduroam.chalmers.se.60379