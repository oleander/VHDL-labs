linus@dhcp-074127.eduroam.chalmers.se.43552