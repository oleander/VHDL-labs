linus@linus-oleanders-macbook.local.980