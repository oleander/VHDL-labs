linus@dhcp-076097.eduroam.chalmers.se.35440