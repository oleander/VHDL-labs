linus@linus-oleanders-macbook.local.791