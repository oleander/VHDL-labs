linus@dhcp-079030.eduroam.chalmers.se.9922