linus@banan.olf.sgsnet.se.4195