linus@linus-oleanders-macbook.local.17339