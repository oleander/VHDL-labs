linus@dhcp-079070.eduroam.chalmers.se.41930