linus@linus-oleanders-macbook.local.16289