linus@linus-oleanders-macbook.local.18289