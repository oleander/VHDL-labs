linus@dhcp-075075.eduroam.chalmers.se.6746