linus@dhcp-075075.eduroam.chalmers.se.8928