linus@dhcp-074169.eduroam.chalmers.se.69458