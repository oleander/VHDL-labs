linus@dhcp-075075.eduroam.chalmers.se.2144