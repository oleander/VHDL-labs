linus@linus-oleanders-macbook.local.3672