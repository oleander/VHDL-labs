linus@dhcp-075015.eduroam.chalmers.se.23945